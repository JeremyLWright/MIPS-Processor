`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:15:23 11/11/2007 
// Design Name: 
// Module Name:    ShiftLeft2_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ShiftLeft2_tb();

reg [31:0] a_t;
wire [31:0] result_t;

//ShiftLeft2 ShiftLeft2_t(a_t, result_t);

initial 
	begin 
		a_t <= 1;
		
	end
	


endmodule
