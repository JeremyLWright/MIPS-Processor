`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:38:43 11/10/2007 
// Design Name: 
// Module Name:    ANDGate_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ANDGate_tb();

reg a_t,b_t;
wire result_t;

//ANDGate ANDGate1(a_t, b_t, result_t);

initial 
	begin 
		a_t <= 0;
		b_t <= 0;
	end

endmodule
