`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:40:10 10/13/2007 
// Design Name: 
// Module Name:    DataMemory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DataMemory(Address, WriteData, MemRead, MemWrite, Clk, ReadData);

input [31:0] Address; // 32-bit address to memory.
input [31:0] WriteData; // Data to be written into WriteRegister
input MemRead; // Data in memory location Address is read if
					// this control is set

input Clk;
input MemWrite; // WriteData is written in Address during
					// positive clock edge if this control is set
					
output [31:0] ReadData; // Value read from memory location Address

reg [31:0] ReadData;  //output register 

//data memory registers for storage. reg initialization ends at line 518
reg [31:0] dm000, dm001, dm002, dm003, dm004, dm005, dm006, dm007, dm008, dm009, dm010,
			  dm011, dm012, dm013, dm014, dm015, dm016, dm017, dm018, dm019, dm020, dm021,
			  dm022, dm023, dm024, dm025, dm026, dm027, dm028, dm029, dm030, dm031, dm032,
				dm033, dm034, dm035, dm036, dm037, dm038, dm039, dm040, dm041, dm042, dm043,
				dm044, dm045, dm046, dm047, dm048, dm049, dm050, dm051, dm052, dm053, dm054,
				dm055, dm056, dm057, dm058, dm059, dm060, dm061,
dm062,
dm063,
dm064,
dm065,
dm066,
dm067,
dm068,
dm069,
dm070,
dm071,
dm072,
dm073,
dm074,
dm075,
dm076,
dm077,
dm078,
dm079,
dm080,
dm081,
dm082,
dm083,
dm084,
dm085,
dm086,
dm087,
dm088,
dm089,
dm090,
dm091,
dm092,
dm093,
dm094,
dm095,
dm096,
dm097,
dm098,
dm099,
dm100,
dm101,
dm102,
dm103,
dm104,
dm105,
dm106,
dm107,
dm108,
dm109,
dm110,
dm111,
dm112,
dm113,
dm114,
dm115,
dm116,
dm117,
dm118,
dm119,
dm120,
dm121,
dm122,
dm123,
dm124,
dm125,
dm126,
dm127,
dm128,
dm129,
dm130,
dm131,
dm132,
dm133,
dm134,
dm135,
dm136,
dm137,
dm138,
dm139,
dm140,
dm141,
dm142,
dm143,
dm144,
dm145,
dm146,
dm147,
dm148,
dm149,
dm150,
dm151,
dm152,
dm153,
dm154,
dm155,
dm156,
dm157,
dm158,
dm159,
dm160,
dm161,
dm162,
dm163,
dm164,
dm165,
dm166,
dm167,
dm168,
dm169,
dm170,
dm171,
dm172,
dm173,
dm174,
dm175,
dm176,
dm177,
dm178,
dm179,
dm180,
dm181,
dm182,
dm183,
dm184,
dm185,
dm186,
dm187,
dm188,
dm189,
dm190,
dm191,
dm192,
dm193,
dm194,
dm195,
dm196,
dm197,
dm198,
dm199,
dm200,
dm201,
dm202,
dm203,
dm204,
dm205,
dm206,
dm207,
dm208,
dm209,
dm210,
dm211,
dm212,
dm213,
dm214,
dm215,
dm216,
dm217,
dm218,
dm219,
dm220,
dm221,
dm222,
dm223,
dm224,
dm225,
dm226,
dm227,
dm228,
dm229,
dm230,
dm231,
dm232,
dm233,
dm234,
dm235,
dm236,
dm237,
dm238,
dm239,
dm240,
dm241,
dm242,
dm243,
dm244,
dm245,
dm246,
dm247,
dm248,
dm249,
dm250,
dm251,
dm252,
dm253,
dm254,
dm255,
dm256,
dm257,
dm258,
dm259,
dm260,
dm261,
dm262,
dm263,
dm264,
dm265,
dm266,
dm267,
dm268,
dm269,
dm270,
dm271,
dm272,
dm273,
dm274,
dm275,
dm276,
dm277,
dm278,
dm279,
dm280,
dm281,
dm282,
dm283,
dm284,
dm285,
dm286,
dm287,
dm288,
dm289,
dm290,
dm291,
dm292,
dm293,
dm294,
dm295,
dm296,
dm297,
dm298,
dm299,
dm300,
dm301,
dm302,
dm303,
dm304,
dm305,
dm306,
dm307,
dm308,
dm309,
dm310,
dm311,
dm312,
dm313,
dm314,
dm315,
dm316,
dm317,
dm318,
dm319,
dm320,
dm321,
dm322,
dm323,
dm324,
dm325,
dm326,
dm327,
dm328,
dm329,
dm330,
dm331,
dm332,
dm333,
dm334,
dm335,
dm336,
dm337,
dm338,
dm339,
dm340,
dm341,
dm342,
dm343,
dm344,
dm345,
dm346,
dm347,
dm348,
dm349,
dm350,
dm351,
dm352,
dm353,
dm354,
dm355,
dm356,
dm357,
dm358,
dm359,
dm360,
dm361,
dm362,
dm363,
dm364,
dm365,
dm366,
dm367,
dm368,
dm369,
dm370,
dm371,
dm372,
dm373,
dm374,
dm375,
dm376,
dm377,
dm378,
dm379,
dm380,
dm381,
dm382,
dm383,
dm384,
dm385,
dm386,
dm387,
dm388,
dm389,
dm390,
dm391,
dm392,
dm393,
dm394,
dm395,
dm396,
dm397,
dm398,
dm399,
dm400,
dm401,
dm402,
dm403,
dm404,
dm405,
dm406,
dm407,
dm408,
dm409,
dm410,
dm411,
dm412,
dm413,
dm414,
dm415,
dm416,
dm417,
dm418,
dm419,
dm420,
dm421,
dm422,
dm423,
dm424,
dm425,
dm426,
dm427,
dm428,
dm429,
dm430,
dm431,
dm432,
dm433,
dm434,
dm435,
dm436,
dm437,
dm438,
dm439,
dm440,
dm441,
dm442,
dm443,
dm444,
dm445,
dm446,
dm447,
dm448,
dm449,
dm450,
dm451,
dm452,
dm453,
dm454,
dm455,
dm456,
dm457,
dm458,
dm459,
dm460,
dm461,
dm462,
dm463,
dm464,
dm465,
dm466,
dm467,
dm468,
dm469,
dm470,
dm471,
dm472,
dm473,
dm474,
dm475,
dm476,
dm477,
dm478,
dm479,
dm480,
dm481,
dm482,
dm483,
dm484,
dm485,
dm486,
dm487,
dm488,
dm489,
dm490,
dm491,
dm492,
dm493,
dm494,
dm495,
dm496,
dm497,
dm498,
dm499,
dm500,
dm501,
dm502,
dm503,
dm504,
dm505,
dm506,
dm507,
dm508,
dm509,
dm510,
dm511;


initial
	begin
		  dm009 <= 32'b00000000000100011000000000000001;
		  //dm017 <= 32'b00000000000000000000000000000011;
		  //R09 <= 32'b00000010001010010111000000000000;
	end


//always  @ (posedge Clk)// Select mem address and write to that address
always  @ (WriteData or Address)// Select mem address and write to that address

   begin
      if(MemWrite == 1)
			case(Address)   //stops at line 
9'd0: dm000 = WriteData;
9'd1: dm001 = WriteData;
9'd2: dm002 = WriteData;
9'd3: dm003 = WriteData;
9'd4: dm004 = WriteData;
9'd5: dm005 = WriteData;
9'd6: dm006 = WriteData;
9'd7: dm007 = WriteData;
9'd8: dm008 = WriteData;
9'd9: dm009 = WriteData;
9'd10: dm010 = WriteData;
9'd11: dm011 = WriteData;
9'd12: dm012 = WriteData;
9'd13: dm013 = WriteData;
9'd14: dm014 = WriteData;
9'd15: dm015 = WriteData;
9'd16: dm016 = WriteData;
9'd17: dm017 = WriteData;
9'd18: dm018 = WriteData;
9'd19: dm019 = WriteData;
9'd20: dm020 = WriteData;
9'd21: dm021 = WriteData;
9'd22: dm022 = WriteData;
9'd23: dm023 = WriteData;
9'd24: dm024 = WriteData;
9'd25: dm025 = WriteData;
9'd26: dm026 = WriteData;
9'd27: dm027 = WriteData;
9'd28: dm028 = WriteData;
9'd29: dm029 = WriteData;
9'd30: dm030 = WriteData;
9'd31: dm031 = WriteData;
9'd32: dm032 = WriteData;
9'd33: dm033 = WriteData;
9'd34: dm034 = WriteData;
9'd35: dm035 = WriteData;
9'd36: dm036 = WriteData;
9'd37: dm037 = WriteData;
9'd38: dm038 = WriteData;
9'd39: dm039 = WriteData;
9'd40: dm040 = WriteData;
9'd41: dm041 = WriteData;
9'd42: dm042 = WriteData;
9'd43: dm043 = WriteData;
9'd44: dm044 = WriteData;
9'd45: dm045 = WriteData;
9'd46: dm046 = WriteData;
9'd47: dm047 = WriteData;
9'd48: dm048 = WriteData;
9'd49: dm049 = WriteData;
9'd50: dm050 = WriteData;
9'd51: dm051 = WriteData;
9'd52: dm052 = WriteData;
9'd53: dm053 = WriteData;
9'd54: dm054 = WriteData;
9'd55: dm055 = WriteData;
9'd56: dm056 = WriteData;
9'd57: dm057 = WriteData;
9'd58: dm058 = WriteData;
9'd59: dm059 = WriteData;
9'd60: dm060 = WriteData;
9'd61: dm061 = WriteData;
9'd62: dm062 = WriteData;
9'd63: dm063 = WriteData;
9'd64: dm064 = WriteData;
9'd65: dm065 = WriteData;
9'd66: dm066 = WriteData;
9'd67: dm067 = WriteData;
9'd68: dm068 = WriteData;
9'd69: dm069 = WriteData;
9'd70: dm070 = WriteData;
9'd71: dm071 = WriteData;
9'd72: dm072 = WriteData;
9'd73: dm073 = WriteData;
9'd74: dm074 = WriteData;
9'd75: dm075 = WriteData;
9'd76: dm076 = WriteData;
9'd77: dm077 = WriteData;
9'd78: dm078 = WriteData;
9'd79: dm079 = WriteData;
9'd80: dm080 = WriteData;
9'd81: dm081 = WriteData;
9'd82: dm082 = WriteData;
9'd83: dm083 = WriteData;
9'd84: dm084 = WriteData;
9'd85: dm085 = WriteData;
9'd86: dm086 = WriteData;
9'd87: dm087 = WriteData;
9'd88: dm088 = WriteData;
9'd89: dm089 = WriteData;
9'd90: dm090 = WriteData;
9'd91: dm091 = WriteData;
9'd92: dm092 = WriteData;
9'd93: dm093 = WriteData;
9'd94: dm094 = WriteData;
9'd95: dm095 = WriteData;
9'd96: dm096 = WriteData;
9'd97: dm097 = WriteData;
9'd98: dm098 = WriteData;
9'd99: dm099 = WriteData;
9'd100: dm100 = WriteData;
9'd101: dm101 = WriteData;
9'd102: dm102 = WriteData;
9'd103: dm103 = WriteData;
9'd104: dm104 = WriteData;
9'd105: dm105 = WriteData;
9'd106: dm106 = WriteData;
9'd107: dm107 = WriteData;
9'd108: dm108 = WriteData;
9'd109: dm109 = WriteData;
9'd110: dm110 = WriteData;
9'd111: dm111 = WriteData;
9'd112: dm112 = WriteData;
9'd113: dm113 = WriteData;
9'd114: dm114 = WriteData;
9'd115: dm115 = WriteData;
9'd116: dm116 = WriteData;
9'd117: dm117 = WriteData;
9'd118: dm118 = WriteData;
9'd119: dm119 = WriteData;
9'd120: dm120 = WriteData;
9'd121: dm121 = WriteData;
9'd122: dm122 = WriteData;
9'd123: dm123 = WriteData;
9'd124: dm124 = WriteData;
9'd125: dm125 = WriteData;
9'd126: dm126 = WriteData;
9'd127: dm127 = WriteData;
9'd128: dm128 = WriteData;
9'd129: dm129 = WriteData;
9'd130: dm130 = WriteData;
9'd131: dm131 = WriteData;
9'd132: dm132 = WriteData;
9'd133: dm133 = WriteData;
9'd134: dm134 = WriteData;
9'd135: dm135 = WriteData;
9'd136: dm136 = WriteData;
9'd137: dm137 = WriteData;
9'd138: dm138 = WriteData;
9'd139: dm139 = WriteData;
9'd140: dm140 = WriteData;
9'd141: dm141 = WriteData;
9'd142: dm142 = WriteData;
9'd143: dm143 = WriteData;
9'd144: dm144 = WriteData;
9'd145: dm145 = WriteData;
9'd146: dm146 = WriteData;
9'd147: dm147 = WriteData;
9'd148: dm148 = WriteData;
9'd149: dm149 = WriteData;
9'd150: dm150 = WriteData;
9'd151: dm151 = WriteData;
9'd152: dm152 = WriteData;
9'd153: dm153 = WriteData;
9'd154: dm154 = WriteData;
9'd155: dm155 = WriteData;
9'd156: dm156 = WriteData;
9'd157: dm157 = WriteData;
9'd158: dm158 = WriteData;
9'd159: dm159 = WriteData;
9'd160: dm160 = WriteData;
9'd161: dm161 = WriteData;
9'd162: dm162 = WriteData;
9'd163: dm163 = WriteData;
9'd164: dm164 = WriteData;
9'd165: dm165 = WriteData;
9'd166: dm166 = WriteData;
9'd167: dm167 = WriteData;
9'd168: dm168 = WriteData;
9'd169: dm169 = WriteData;
9'd170: dm170 = WriteData;
9'd171: dm171 = WriteData;
9'd172: dm172 = WriteData;
9'd173: dm173 = WriteData;
9'd174: dm174 = WriteData;
9'd175: dm175 = WriteData;
9'd176: dm176 = WriteData;
9'd177: dm177 = WriteData;
9'd178: dm178 = WriteData;
9'd179: dm179 = WriteData;
9'd180: dm180 = WriteData;
9'd181: dm181 = WriteData;
9'd182: dm182 = WriteData;
9'd183: dm183 = WriteData;
9'd184: dm184 = WriteData;
9'd185: dm185 = WriteData;
9'd186: dm186 = WriteData;
9'd187: dm187 = WriteData;
9'd188: dm188 = WriteData;
9'd189: dm189 = WriteData;
9'd190: dm190 = WriteData;
9'd191: dm191 = WriteData;
9'd192: dm192 = WriteData;
9'd193: dm193 = WriteData;
9'd194: dm194 = WriteData;
9'd195: dm195 = WriteData;
9'd196: dm196 = WriteData;
9'd197: dm197 = WriteData;
9'd198: dm198 = WriteData;
9'd199: dm199 = WriteData;
9'd200: dm200 = WriteData;
9'd201: dm201 = WriteData;
9'd202: dm202 = WriteData;
9'd203: dm203 = WriteData;
9'd204: dm204 = WriteData;
9'd205: dm205 = WriteData;
9'd206: dm206 = WriteData;
9'd207: dm207 = WriteData;
9'd208: dm208 = WriteData;
9'd209: dm209 = WriteData;
9'd210: dm210 = WriteData;
9'd211: dm211 = WriteData;
9'd212: dm212 = WriteData;
9'd213: dm213 = WriteData;
9'd214: dm214 = WriteData;
9'd215: dm215 = WriteData;
9'd216: dm216 = WriteData;
9'd217: dm217 = WriteData;
9'd218: dm218 = WriteData;
9'd219: dm219 = WriteData;
9'd220: dm220 = WriteData;
9'd221: dm221 = WriteData;
9'd222: dm222 = WriteData;
9'd223: dm223 = WriteData;
9'd224: dm224 = WriteData;
9'd225: dm225 = WriteData;
9'd226: dm226 = WriteData;
9'd227: dm227 = WriteData;
9'd228: dm228 = WriteData;
9'd229: dm229 = WriteData;
9'd230: dm230 = WriteData;
9'd231: dm231 = WriteData;
9'd232: dm232 = WriteData;
9'd233: dm233 = WriteData;
9'd234: dm234 = WriteData;
9'd235: dm235 = WriteData;
9'd236: dm236 = WriteData;
9'd237: dm237 = WriteData;
9'd238: dm238 = WriteData;
9'd239: dm239 = WriteData;
9'd240: dm240 = WriteData;
9'd241: dm241 = WriteData;
9'd242: dm242 = WriteData;
9'd243: dm243 = WriteData;
9'd244: dm244 = WriteData;
9'd245: dm245 = WriteData;
9'd246: dm246 = WriteData;
9'd247: dm247 = WriteData;
9'd248: dm248 = WriteData;
9'd249: dm249 = WriteData;
9'd250: dm250 = WriteData;
9'd251: dm251 = WriteData;
9'd252: dm252 = WriteData;
9'd253: dm253 = WriteData;
9'd254: dm254 = WriteData;
9'd255: dm255 = WriteData;
9'd256: dm256 = WriteData;
9'd257: dm257 = WriteData;
9'd258: dm258 = WriteData;
9'd259: dm259 = WriteData;
9'd260: dm260 = WriteData;
9'd261: dm261 = WriteData;
9'd262: dm262 = WriteData;
9'd263: dm263 = WriteData;
9'd264: dm264 = WriteData;
9'd265: dm265 = WriteData;
9'd266: dm266 = WriteData;
9'd267: dm267 = WriteData;
9'd268: dm268 = WriteData;
9'd269: dm269 = WriteData;
9'd270: dm270 = WriteData;
9'd271: dm271 = WriteData;
9'd272: dm272 = WriteData;
9'd273: dm273 = WriteData;
9'd274: dm274 = WriteData;
9'd275: dm275 = WriteData;
9'd276: dm276 = WriteData;
9'd277: dm277 = WriteData;
9'd278: dm278 = WriteData;
9'd279: dm279 = WriteData;
9'd280: dm280 = WriteData;
9'd281: dm281 = WriteData;
9'd282: dm282 = WriteData;
9'd283: dm283 = WriteData;
9'd284: dm284 = WriteData;
9'd285: dm285 = WriteData;
9'd286: dm286 = WriteData;
9'd287: dm287 = WriteData;
9'd288: dm288 = WriteData;
9'd289: dm289 = WriteData;
9'd290: dm290 = WriteData;
9'd291: dm291 = WriteData;
9'd292: dm292 = WriteData;
9'd293: dm293 = WriteData;
9'd294: dm294 = WriteData;
9'd295: dm295 = WriteData;
9'd296: dm296 = WriteData;
9'd297: dm297 = WriteData;
9'd298: dm298 = WriteData;
9'd299: dm299 = WriteData;
9'd300: dm300 = WriteData;
9'd301: dm301 = WriteData;
9'd302: dm302 = WriteData;
9'd303: dm303 = WriteData;
9'd304: dm304 = WriteData;
9'd305: dm305 = WriteData;
9'd306: dm306 = WriteData;
9'd307: dm307 = WriteData;
9'd308: dm308 = WriteData;
9'd309: dm309 = WriteData;
9'd310: dm310 = WriteData;
9'd311: dm311 = WriteData;
9'd312: dm312 = WriteData;
9'd313: dm313 = WriteData;
9'd314: dm314 = WriteData;
9'd315: dm315 = WriteData;
9'd316: dm316 = WriteData;
9'd317: dm317 = WriteData;
9'd318: dm318 = WriteData;
9'd319: dm319 = WriteData;
9'd320: dm320 = WriteData;
9'd321: dm321 = WriteData;
9'd322: dm322 = WriteData;
9'd323: dm323 = WriteData;
9'd324: dm324 = WriteData;
9'd325: dm325 = WriteData;
9'd326: dm326 = WriteData;
9'd327: dm327 = WriteData;
9'd328: dm328 = WriteData;
9'd329: dm329 = WriteData;
9'd330: dm330 = WriteData;
9'd331: dm331 = WriteData;
9'd332: dm332 = WriteData;
9'd333: dm333 = WriteData;
9'd334: dm334 = WriteData;
9'd335: dm335 = WriteData;
9'd336: dm336 = WriteData;
9'd337: dm337 = WriteData;
9'd338: dm338 = WriteData;
9'd339: dm339 = WriteData;
9'd340: dm340 = WriteData;
9'd341: dm341 = WriteData;
9'd342: dm342 = WriteData;
9'd343: dm343 = WriteData;
9'd344: dm344 = WriteData;
9'd345: dm345 = WriteData;
9'd346: dm346 = WriteData;
9'd347: dm347 = WriteData;
9'd348: dm348 = WriteData;
9'd349: dm349 = WriteData;
9'd350: dm350 = WriteData;
9'd351: dm351 = WriteData;
9'd352: dm352 = WriteData;
9'd353: dm353 = WriteData;
9'd354: dm354 = WriteData;
9'd355: dm355 = WriteData;
9'd356: dm356 = WriteData;
9'd357: dm357 = WriteData;
9'd358: dm358 = WriteData;
9'd359: dm359 = WriteData;
9'd360: dm360 = WriteData;
9'd361: dm361 = WriteData;
9'd362: dm362 = WriteData;
9'd363: dm363 = WriteData;
9'd364: dm364 = WriteData;
9'd365: dm365 = WriteData;
9'd366: dm366 = WriteData;
9'd367: dm367 = WriteData;
9'd368: dm368 = WriteData;
9'd369: dm369 = WriteData;
9'd370: dm370 = WriteData;
9'd371: dm371 = WriteData;
9'd372: dm372 = WriteData;
9'd373: dm373 = WriteData;
9'd374: dm374 = WriteData;
9'd375: dm375 = WriteData;
9'd376: dm376 = WriteData;
9'd377: dm377 = WriteData;
9'd378: dm378 = WriteData;
9'd379: dm379 = WriteData;
9'd380: dm380 = WriteData;
9'd381: dm381 = WriteData;
9'd382: dm382 = WriteData;
9'd383: dm383 = WriteData;
9'd384: dm384 = WriteData;
9'd385: dm385 = WriteData;
9'd386: dm386 = WriteData;
9'd387: dm387 = WriteData;
9'd388: dm388 = WriteData;
9'd389: dm389 = WriteData;
9'd390: dm390 = WriteData;
9'd391: dm391 = WriteData;
9'd392: dm392 = WriteData;
9'd393: dm393 = WriteData;
9'd394: dm394 = WriteData;
9'd395: dm395 = WriteData;
9'd396: dm396 = WriteData;
9'd397: dm397 = WriteData;
9'd398: dm398 = WriteData;
9'd399: dm399 = WriteData;
9'd400: dm400 = WriteData;
9'd401: dm401 = WriteData;
9'd402: dm402 = WriteData;
9'd403: dm403 = WriteData;
9'd404: dm404 = WriteData;
9'd405: dm405 = WriteData;
9'd406: dm406 = WriteData;
9'd407: dm407 = WriteData;
9'd408: dm408 = WriteData;
9'd409: dm409 = WriteData;
9'd410: dm410 = WriteData;
9'd411: dm411 = WriteData;
9'd412: dm412 = WriteData;
9'd413: dm413 = WriteData;
9'd414: dm414 = WriteData;
9'd415: dm415 = WriteData;
9'd416: dm416 = WriteData;
9'd417: dm417 = WriteData;
9'd418: dm418 = WriteData;
9'd419: dm419 = WriteData;
9'd420: dm420 = WriteData;
9'd421: dm421 = WriteData;
9'd422: dm422 = WriteData;
9'd423: dm423 = WriteData;
9'd424: dm424 = WriteData;
9'd425: dm425 = WriteData;
9'd426: dm426 = WriteData;
9'd427: dm427 = WriteData;
9'd428: dm428 = WriteData;
9'd429: dm429 = WriteData;
9'd430: dm430 = WriteData;
9'd431: dm431 = WriteData;
9'd432: dm432 = WriteData;
9'd433: dm433 = WriteData;
9'd434: dm434 = WriteData;
9'd435: dm435 = WriteData;
9'd436: dm436 = WriteData;
9'd437: dm437 = WriteData;
9'd438: dm438 = WriteData;
9'd439: dm439 = WriteData;
9'd440: dm440 = WriteData;
9'd441: dm441 = WriteData;
9'd442: dm442 = WriteData;
9'd443: dm443 = WriteData;
9'd444: dm444 = WriteData;
9'd445: dm445 = WriteData;
9'd446: dm446 = WriteData;
9'd447: dm447 = WriteData;
9'd448: dm448 = WriteData;
9'd449: dm449 = WriteData;
9'd450: dm450 = WriteData;
9'd451: dm451 = WriteData;
9'd452: dm452 = WriteData;
9'd453: dm453 = WriteData;
9'd454: dm454 = WriteData;
9'd455: dm455 = WriteData;
9'd456: dm456 = WriteData;
9'd457: dm457 = WriteData;
9'd458: dm458 = WriteData;
9'd459: dm459 = WriteData;
9'd460: dm460 = WriteData;
9'd461: dm461 = WriteData;
9'd462: dm462 = WriteData;
9'd463: dm463 = WriteData;
9'd464: dm464 = WriteData;
9'd465: dm465 = WriteData;
9'd466: dm466 = WriteData;
9'd467: dm467 = WriteData;
9'd468: dm468 = WriteData;
9'd469: dm469 = WriteData;
9'd470: dm470 = WriteData;
9'd471: dm471 = WriteData;
9'd472: dm472 = WriteData;
9'd473: dm473 = WriteData;
9'd474: dm474 = WriteData;
9'd475: dm475 = WriteData;
9'd476: dm476 = WriteData;
9'd477: dm477 = WriteData;
9'd478: dm478 = WriteData;
9'd479: dm479 = WriteData;
9'd480: dm480 = WriteData;
9'd481: dm481 = WriteData;
9'd482: dm482 = WriteData;
9'd483: dm483 = WriteData;
9'd484: dm484 = WriteData;
9'd485: dm485 = WriteData;
9'd486: dm486 = WriteData;
9'd487: dm487 = WriteData;
9'd488: dm488 = WriteData;
9'd489: dm489 = WriteData;
9'd490: dm490 = WriteData;
9'd491: dm491 = WriteData;
9'd492: dm492 = WriteData;
9'd493: dm493 = WriteData;
9'd494: dm494 = WriteData;
9'd495: dm495 = WriteData;
9'd496: dm496 = WriteData;
9'd497: dm497 = WriteData;
9'd498: dm498 = WriteData;
9'd499: dm499 = WriteData;
9'd500: dm500 = WriteData;
9'd501: dm501 = WriteData;
9'd502: dm502 = WriteData;
9'd503: dm503 = WriteData;
9'd504: dm504 = WriteData;
9'd505: dm505 = WriteData;
9'd506: dm506 = WriteData;
9'd507: dm507 = WriteData;
9'd508: dm508 = WriteData;
9'd509: dm509 = WriteData;
9'd510: dm510 = WriteData;
9'd511: dm511 = WriteData;
endcase
end


//always  @ (negedge Clk)// Select mem space and output on readdata
always  @ (Address)
   begin
      if(MemRead == 1)
			case(Address)   //stops at line 1554
9'd0: ReadData  = dm000;
9'd1: ReadData  = dm001;
9'd2: ReadData  = dm002;
9'd3: ReadData  = dm003;
9'd4: ReadData  = dm004;
9'd5: ReadData  = dm005;
9'd6: ReadData  = dm006;
9'd7: ReadData  = dm007;
9'd8: ReadData  = dm008;
9'd9: ReadData  = dm009;
9'd10: ReadData  = dm010;
9'd11: ReadData  = dm011;
9'd12: ReadData  = dm012;
9'd13: ReadData  = dm013;
9'd14: ReadData  = dm014;
9'd15: ReadData  = dm015;
9'd16: ReadData  = dm016;
9'd17: ReadData  = dm017;
9'd18: ReadData  = dm018;
9'd19: ReadData  = dm019;
9'd20: ReadData  = dm020;
9'd21: ReadData  = dm021;
9'd22: ReadData  = dm022;
9'd23: ReadData  = dm023;
9'd24: ReadData  = dm024;
9'd25: ReadData  = dm025;
9'd26: ReadData  = dm026;
9'd27: ReadData  = dm027;
9'd28: ReadData  = dm028;
9'd29: ReadData  = dm029;
9'd30: ReadData  = dm030;
9'd31: ReadData  = dm031;
9'd32: ReadData  = dm032;
9'd33: ReadData  = dm033;
9'd34: ReadData  = dm034;
9'd35: ReadData  = dm035;
9'd36: ReadData  = dm036;
9'd37: ReadData  = dm037;
9'd38: ReadData  = dm038;
9'd39: ReadData  = dm039;
9'd40: ReadData  = dm040;
9'd41: ReadData  = dm041;
9'd42: ReadData  = dm042;
9'd43: ReadData  = dm043;
9'd44: ReadData  = dm044;
9'd45: ReadData  = dm045;
9'd46: ReadData  = dm046;
9'd47: ReadData  = dm047;
9'd48: ReadData  = dm048;
9'd49: ReadData  = dm049;
9'd50: ReadData  = dm050;
9'd51: ReadData  = dm051;
9'd52: ReadData  = dm052;
9'd53: ReadData  = dm053;
9'd54: ReadData  = dm054;
9'd55: ReadData  = dm055;
9'd56: ReadData  = dm056;
9'd57: ReadData  = dm057;
9'd58: ReadData  = dm058;
9'd59: ReadData  = dm059;
9'd60: ReadData  = dm060;
9'd61: ReadData  = dm061;
9'd62: ReadData  = dm062;
9'd63: ReadData  = dm063;
9'd64: ReadData  = dm064;
9'd65: ReadData  = dm065;
9'd66: ReadData  = dm066;
9'd67: ReadData  = dm067;
9'd68: ReadData  = dm068;
9'd69: ReadData  = dm069;
9'd70: ReadData  = dm070;
9'd71: ReadData  = dm071;
9'd72: ReadData  = dm072;
9'd73: ReadData  = dm073;
9'd74: ReadData  = dm074;
9'd75: ReadData  = dm075;
9'd76: ReadData  = dm076;
9'd77: ReadData  = dm077;
9'd78: ReadData  = dm078;
9'd79: ReadData  = dm079;
9'd80: ReadData  = dm080;
9'd81: ReadData  = dm081;
9'd82: ReadData  = dm082;
9'd83: ReadData  = dm083;
9'd84: ReadData  = dm084;
9'd85: ReadData  = dm085;
9'd86: ReadData  = dm086;
9'd87: ReadData  = dm087;
9'd88: ReadData  = dm088;
9'd89: ReadData  = dm089;
9'd90: ReadData  = dm090;
9'd91: ReadData  = dm091;
9'd92: ReadData  = dm092;
9'd93: ReadData  = dm093;
9'd94: ReadData  = dm094;
9'd95: ReadData  = dm095;
9'd96: ReadData  = dm096;
9'd97: ReadData  = dm097;
9'd98: ReadData  = dm098;
9'd99: ReadData  = dm099;
9'd100: ReadData  = dm100;
9'd101: ReadData  = dm101;
9'd102: ReadData  = dm102;
9'd103: ReadData  = dm103;
9'd104: ReadData  = dm104;
9'd105: ReadData  = dm105;
9'd106: ReadData  = dm106;
9'd107: ReadData  = dm107;
9'd108: ReadData  = dm108;
9'd109: ReadData  = dm109;
9'd110: ReadData  = dm110;
9'd111: ReadData  = dm111;
9'd112: ReadData  = dm112;
9'd113: ReadData  = dm113;
9'd114: ReadData  = dm114;
9'd115: ReadData  = dm115;
9'd116: ReadData  = dm116;
9'd117: ReadData  = dm117;
9'd118: ReadData  = dm118;
9'd119: ReadData  = dm119;
9'd120: ReadData  = dm120;
9'd121: ReadData  = dm121;
9'd122: ReadData  = dm122;
9'd123: ReadData  = dm123;
9'd124: ReadData  = dm124;
9'd125: ReadData  = dm125;
9'd126: ReadData  = dm126;
9'd127: ReadData  = dm127;
9'd128: ReadData  = dm128;
9'd129: ReadData  = dm129;
9'd130: ReadData  = dm130;
9'd131: ReadData  = dm131;
9'd132: ReadData  = dm132;
9'd133: ReadData  = dm133;
9'd134: ReadData  = dm134;
9'd135: ReadData  = dm135;
9'd136: ReadData  = dm136;
9'd137: ReadData  = dm137;
9'd138: ReadData  = dm138;
9'd139: ReadData  = dm139;
9'd140: ReadData  = dm140;
9'd141: ReadData  = dm141;
9'd142: ReadData  = dm142;
9'd143: ReadData  = dm143;
9'd144: ReadData  = dm144;
9'd145: ReadData  = dm145;
9'd146: ReadData  = dm146;
9'd147: ReadData  = dm147;
9'd148: ReadData  = dm148;
9'd149: ReadData  = dm149;
9'd150: ReadData  = dm150;
9'd151: ReadData  = dm151;
9'd152: ReadData  = dm152;
9'd153: ReadData  = dm153;
9'd154: ReadData  = dm154;
9'd155: ReadData  = dm155;
9'd156: ReadData  = dm156;
9'd157: ReadData  = dm157;
9'd158: ReadData  = dm158;
9'd159: ReadData  = dm159;
9'd160: ReadData  = dm160;
9'd161: ReadData  = dm161;
9'd162: ReadData  = dm162;
9'd163: ReadData  = dm163;
9'd164: ReadData  = dm164;
9'd165: ReadData  = dm165;
9'd166: ReadData  = dm166;
9'd167: ReadData  = dm167;
9'd168: ReadData  = dm168;
9'd169: ReadData  = dm169;
9'd170: ReadData  = dm170;
9'd171: ReadData  = dm171;
9'd172: ReadData  = dm172;
9'd173: ReadData  = dm173;
9'd174: ReadData  = dm174;
9'd175: ReadData  = dm175;
9'd176: ReadData  = dm176;
9'd177: ReadData  = dm177;
9'd178: ReadData  = dm178;
9'd179: ReadData  = dm179;
9'd180: ReadData  = dm180;
9'd181: ReadData  = dm181;
9'd182: ReadData  = dm182;
9'd183: ReadData  = dm183;
9'd184: ReadData  = dm184;
9'd185: ReadData  = dm185;
9'd186: ReadData  = dm186;
9'd187: ReadData  = dm187;
9'd188: ReadData  = dm188;
9'd189: ReadData  = dm189;
9'd190: ReadData  = dm190;
9'd191: ReadData  = dm191;
9'd192: ReadData  = dm192;
9'd193: ReadData  = dm193;
9'd194: ReadData  = dm194;
9'd195: ReadData  = dm195;
9'd196: ReadData  = dm196;
9'd197: ReadData  = dm197;
9'd198: ReadData  = dm198;
9'd199: ReadData  = dm199;
9'd200: ReadData  = dm200;
9'd201: ReadData  = dm201;
9'd202: ReadData  = dm202;
9'd203: ReadData  = dm203;
9'd204: ReadData  = dm204;
9'd205: ReadData  = dm205;
9'd206: ReadData  = dm206;
9'd207: ReadData  = dm207;
9'd208: ReadData  = dm208;
9'd209: ReadData  = dm209;
9'd210: ReadData  = dm210;
9'd211: ReadData  = dm211;
9'd212: ReadData  = dm212;
9'd213: ReadData  = dm213;
9'd214: ReadData  = dm214;
9'd215: ReadData  = dm215;
9'd216: ReadData  = dm216;
9'd217: ReadData  = dm217;
9'd218: ReadData  = dm218;
9'd219: ReadData  = dm219;
9'd220: ReadData  = dm220;
9'd221: ReadData  = dm221;
9'd222: ReadData  = dm222;
9'd223: ReadData  = dm223;
9'd224: ReadData  = dm224;
9'd225: ReadData  = dm225;
9'd226: ReadData  = dm226;
9'd227: ReadData  = dm227;
9'd228: ReadData  = dm228;
9'd229: ReadData  = dm229;
9'd230: ReadData  = dm230;
9'd231: ReadData  = dm231;
9'd232: ReadData  = dm232;
9'd233: ReadData  = dm233;
9'd234: ReadData  = dm234;
9'd235: ReadData  = dm235;
9'd236: ReadData  = dm236;
9'd237: ReadData  = dm237;
9'd238: ReadData  = dm238;
9'd239: ReadData  = dm239;
9'd240: ReadData  = dm240;
9'd241: ReadData  = dm241;
9'd242: ReadData  = dm242;
9'd243: ReadData  = dm243;
9'd244: ReadData  = dm244;
9'd245: ReadData  = dm245;
9'd246: ReadData  = dm246;
9'd247: ReadData  = dm247;
9'd248: ReadData  = dm248;
9'd249: ReadData  = dm249;
9'd250: ReadData  = dm250;
9'd251: ReadData  = dm251;
9'd252: ReadData  = dm252;
9'd253: ReadData  = dm253;
9'd254: ReadData  = dm254;
9'd255: ReadData  = dm255;
9'd256: ReadData  = dm256;
9'd257: ReadData  = dm257;
9'd258: ReadData  = dm258;
9'd259: ReadData  = dm259;
9'd260: ReadData  = dm260;
9'd261: ReadData  = dm261;
9'd262: ReadData  = dm262;
9'd263: ReadData  = dm263;
9'd264: ReadData  = dm264;
9'd265: ReadData  = dm265;
9'd266: ReadData  = dm266;
9'd267: ReadData  = dm267;
9'd268: ReadData  = dm268;
9'd269: ReadData  = dm269;
9'd270: ReadData  = dm270;
9'd271: ReadData  = dm271;
9'd272: ReadData  = dm272;
9'd273: ReadData  = dm273;
9'd274: ReadData  = dm274;
9'd275: ReadData  = dm275;
9'd276: ReadData  = dm276;
9'd277: ReadData  = dm277;
9'd278: ReadData  = dm278;
9'd279: ReadData  = dm279;
9'd280: ReadData  = dm280;
9'd281: ReadData  = dm281;
9'd282: ReadData  = dm282;
9'd283: ReadData  = dm283;
9'd284: ReadData  = dm284;
9'd285: ReadData  = dm285;
9'd286: ReadData  = dm286;
9'd287: ReadData  = dm287;
9'd288: ReadData  = dm288;
9'd289: ReadData  = dm289;
9'd290: ReadData  = dm290;
9'd291: ReadData  = dm291;
9'd292: ReadData  = dm292;
9'd293: ReadData  = dm293;
9'd294: ReadData  = dm294;
9'd295: ReadData  = dm295;
9'd296: ReadData  = dm296;
9'd297: ReadData  = dm297;
9'd298: ReadData  = dm298;
9'd299: ReadData  = dm299;
9'd300: ReadData  = dm300;
9'd301: ReadData  = dm301;
9'd302: ReadData  = dm302;
9'd303: ReadData  = dm303;
9'd304: ReadData  = dm304;
9'd305: ReadData  = dm305;
9'd306: ReadData  = dm306;
9'd307: ReadData  = dm307;
9'd308: ReadData  = dm308;
9'd309: ReadData  = dm309;
9'd310: ReadData  = dm310;
9'd311: ReadData  = dm311;
9'd312: ReadData  = dm312;
9'd313: ReadData  = dm313;
9'd314: ReadData  = dm314;
9'd315: ReadData  = dm315;
9'd316: ReadData  = dm316;
9'd317: ReadData  = dm317;
9'd318: ReadData  = dm318;
9'd319: ReadData  = dm319;
9'd320: ReadData  = dm320;
9'd321: ReadData  = dm321;
9'd322: ReadData  = dm322;
9'd323: ReadData  = dm323;
9'd324: ReadData  = dm324;
9'd325: ReadData  = dm325;
9'd326: ReadData  = dm326;
9'd327: ReadData  = dm327;
9'd328: ReadData  = dm328;
9'd329: ReadData  = dm329;
9'd330: ReadData  = dm330;
9'd331: ReadData  = dm331;
9'd332: ReadData  = dm332;
9'd333: ReadData  = dm333;
9'd334: ReadData  = dm334;
9'd335: ReadData  = dm335;
9'd336: ReadData  = dm336;
9'd337: ReadData  = dm337;
9'd338: ReadData  = dm338;
9'd339: ReadData  = dm339;
9'd340: ReadData  = dm340;
9'd341: ReadData  = dm341;
9'd342: ReadData  = dm342;
9'd343: ReadData  = dm343;
9'd344: ReadData  = dm344;
9'd345: ReadData  = dm345;
9'd346: ReadData  = dm346;
9'd347: ReadData  = dm347;
9'd348: ReadData  = dm348;
9'd349: ReadData  = dm349;
9'd350: ReadData  = dm350;
9'd351: ReadData  = dm351;
9'd352: ReadData  = dm352;
9'd353: ReadData  = dm353;
9'd354: ReadData  = dm354;
9'd355: ReadData  = dm355;
9'd356: ReadData  = dm356;
9'd357: ReadData  = dm357;
9'd358: ReadData  = dm358;
9'd359: ReadData  = dm359;
9'd360: ReadData  = dm360;
9'd361: ReadData  = dm361;
9'd362: ReadData  = dm362;
9'd363: ReadData  = dm363;
9'd364: ReadData  = dm364;
9'd365: ReadData  = dm365;
9'd366: ReadData  = dm366;
9'd367: ReadData  = dm367;
9'd368: ReadData  = dm368;
9'd369: ReadData  = dm369;
9'd370: ReadData  = dm370;
9'd371: ReadData  = dm371;
9'd372: ReadData  = dm372;
9'd373: ReadData  = dm373;
9'd374: ReadData  = dm374;
9'd375: ReadData  = dm375;
9'd376: ReadData  = dm376;
9'd377: ReadData  = dm377;
9'd378: ReadData  = dm378;
9'd379: ReadData  = dm379;
9'd380: ReadData  = dm380;
9'd381: ReadData  = dm381;
9'd382: ReadData  = dm382;
9'd383: ReadData  = dm383;
9'd384: ReadData  = dm384;
9'd385: ReadData  = dm385;
9'd386: ReadData  = dm386;
9'd387: ReadData  = dm387;
9'd388: ReadData  = dm388;
9'd389: ReadData  = dm389;
9'd390: ReadData  = dm390;
9'd391: ReadData  = dm391;
9'd392: ReadData  = dm392;
9'd393: ReadData  = dm393;
9'd394: ReadData  = dm394;
9'd395: ReadData  = dm395;
9'd396: ReadData  = dm396;
9'd397: ReadData  = dm397;
9'd398: ReadData  = dm398;
9'd399: ReadData  = dm399;
9'd400: ReadData  = dm400;
9'd401: ReadData  = dm401;
9'd402: ReadData  = dm402;
9'd403: ReadData  = dm403;
9'd404: ReadData  = dm404;
9'd405: ReadData  = dm405;
9'd406: ReadData  = dm406;
9'd407: ReadData  = dm407;
9'd408: ReadData  = dm408;
9'd409: ReadData  = dm409;
9'd410: ReadData  = dm410;
9'd411: ReadData  = dm411;
9'd412: ReadData  = dm412;
9'd413: ReadData  = dm413;
9'd414: ReadData  = dm414;
9'd415: ReadData  = dm415;
9'd416: ReadData  = dm416;
9'd417: ReadData  = dm417;
9'd418: ReadData  = dm418;
9'd419: ReadData  = dm419;
9'd420: ReadData  = dm420;
9'd421: ReadData  = dm421;
9'd422: ReadData  = dm422;
9'd423: ReadData  = dm423;
9'd424: ReadData  = dm424;
9'd425: ReadData  = dm425;
9'd426: ReadData  = dm426;
9'd427: ReadData  = dm427;
9'd428: ReadData  = dm428;
9'd429: ReadData  = dm429;
9'd430: ReadData  = dm430;
9'd431: ReadData  = dm431;
9'd432: ReadData  = dm432;
9'd433: ReadData  = dm433;
9'd434: ReadData  = dm434;
9'd435: ReadData  = dm435;
9'd436: ReadData  = dm436;
9'd437: ReadData  = dm437;
9'd438: ReadData  = dm438;
9'd439: ReadData  = dm439;
9'd440: ReadData  = dm440;
9'd441: ReadData  = dm441;
9'd442: ReadData  = dm442;
9'd443: ReadData  = dm443;
9'd444: ReadData  = dm444;
9'd445: ReadData  = dm445;
9'd446: ReadData  = dm446;
9'd447: ReadData  = dm447;
9'd448: ReadData  = dm448;
9'd449: ReadData  = dm449;
9'd450: ReadData  = dm450;
9'd451: ReadData  = dm451;
9'd452: ReadData  = dm452;
9'd453: ReadData  = dm453;
9'd454: ReadData  = dm454;
9'd455: ReadData  = dm455;
9'd456: ReadData  = dm456;
9'd457: ReadData  = dm457;
9'd458: ReadData  = dm458;
9'd459: ReadData  = dm459;
9'd460: ReadData  = dm460;
9'd461: ReadData  = dm461;
9'd462: ReadData  = dm462;
9'd463: ReadData  = dm463;
9'd464: ReadData  = dm464;
9'd465: ReadData  = dm465;
9'd466: ReadData  = dm466;
9'd467: ReadData  = dm467;
9'd468: ReadData  = dm468;
9'd469: ReadData  = dm469;
9'd470: ReadData  = dm470;
9'd471: ReadData  = dm471;
9'd472: ReadData  = dm472;
9'd473: ReadData  = dm473;
9'd474: ReadData  = dm474;
9'd475: ReadData  = dm475;
9'd476: ReadData  = dm476;
9'd477: ReadData  = dm477;
9'd478: ReadData  = dm478;
9'd479: ReadData  = dm479;
9'd480: ReadData  = dm480;
9'd481: ReadData  = dm481;
9'd482: ReadData  = dm482;
9'd483: ReadData  = dm483;
9'd484: ReadData  = dm484;
9'd485: ReadData  = dm485;
9'd486: ReadData  = dm486;
9'd487: ReadData  = dm487;
9'd488: ReadData  = dm488;
9'd489: ReadData  = dm489;
9'd490: ReadData  = dm490;
9'd491: ReadData  = dm491;
9'd492: ReadData  = dm492;
9'd493: ReadData  = dm493;
9'd494: ReadData  = dm494;
9'd495: ReadData  = dm495;
9'd496: ReadData  = dm496;
9'd497: ReadData  = dm497;
9'd498: ReadData  = dm498;
9'd499: ReadData  = dm499;
9'd500: ReadData  = dm500;
9'd501: ReadData  = dm501;
9'd502: ReadData  = dm502;
9'd503: ReadData  = dm503;
9'd504: ReadData  = dm504;
9'd505: ReadData  = dm505;
9'd506: ReadData  = dm506;
9'd507: ReadData  = dm507;
9'd508: ReadData  = dm508;
9'd509: ReadData  = dm509;
9'd510: ReadData  = dm510;
9'd511: ReadData  = dm511;

endcase
end



always @ (MemRead == 0)  // No read or write output 0 on readdata. 
   begin
      if(MemRead == 0)
			case(Address)   //stops at line 
9'd0: ReadData = 0;
9'd1: ReadData = 0;
9'd2: ReadData = 0;
9'd3: ReadData = 0;
9'd4: ReadData = 0;
9'd5: ReadData = 0;
9'd6: ReadData = 0;
9'd7: ReadData = 0;
9'd8: ReadData = 0;
9'd9: ReadData = 0;
9'd10: ReadData = 0;
9'd11: ReadData = 0;
9'd12: ReadData = 0;
9'd13: ReadData = 0;
9'd14: ReadData = 0;
9'd15: ReadData = 0;
9'd16: ReadData = 0;
9'd17: ReadData = 0;
9'd18: ReadData = 0;
9'd19: ReadData = 0;
9'd20: ReadData = 0;
9'd21: ReadData = 0;
9'd22: ReadData = 0;
9'd23: ReadData = 0;
9'd24: ReadData = 0;
9'd25: ReadData = 0;
9'd26: ReadData = 0;
9'd27: ReadData = 0;
9'd28: ReadData = 0;
9'd29: ReadData = 0;
9'd30: ReadData = 0;
9'd31: ReadData = 0;
9'd32: ReadData = 0;
9'd33: ReadData = 0;
9'd34: ReadData = 0;
9'd35: ReadData = 0;
9'd36: ReadData = 0;
9'd37: ReadData = 0;
9'd38: ReadData = 0;
9'd39: ReadData = 0;
9'd40: ReadData = 0;
9'd41: ReadData = 0;
9'd42: ReadData = 0;
9'd43: ReadData = 0;
9'd44: ReadData = 0;
9'd45: ReadData = 0;
9'd46: ReadData = 0;
9'd47: ReadData = 0;
9'd48: ReadData = 0;
9'd49: ReadData = 0;
9'd50: ReadData = 0;
9'd51: ReadData = 0;
9'd52: ReadData = 0;
9'd53: ReadData = 0;
9'd54: ReadData = 0;
9'd55: ReadData = 0;
9'd56: ReadData = 0;
9'd57: ReadData = 0;
9'd58: ReadData = 0;
9'd59: ReadData = 0;
9'd60: ReadData = 0;
9'd61: ReadData = 0;
9'd62: ReadData = 0;
9'd63: ReadData = 0;
9'd64: ReadData = 0;
9'd65: ReadData = 0;
9'd66: ReadData = 0;
9'd67: ReadData = 0;
9'd68: ReadData = 0;
9'd69: ReadData = 0;
9'd70: ReadData = 0;
9'd71: ReadData = 0;
9'd72: ReadData = 0;
9'd73: ReadData = 0;
9'd74: ReadData = 0;
9'd75: ReadData = 0;
9'd76: ReadData = 0;
9'd77: ReadData = 0;
9'd78: ReadData = 0;
9'd79: ReadData = 0;
9'd80: ReadData = 0;
9'd81: ReadData = 0;
9'd82: ReadData = 0;
9'd83: ReadData = 0;
9'd84: ReadData = 0;
9'd85: ReadData = 0;
9'd86: ReadData = 0;
9'd87: ReadData = 0;
9'd88: ReadData = 0;
9'd89: ReadData = 0;
9'd90: ReadData = 0;
9'd91: ReadData = 0;
9'd92: ReadData = 0;
9'd93: ReadData = 0;
9'd94: ReadData = 0;
9'd95: ReadData = 0;
9'd96: ReadData = 0;
9'd97: ReadData = 0;
9'd98: ReadData = 0;
9'd99: ReadData = 0;
9'd100: ReadData = 0;
9'd101: ReadData = 0;
9'd102: ReadData = 0;
9'd103: ReadData = 0;
9'd104: ReadData = 0;
9'd105: ReadData = 0;
9'd106: ReadData = 0;
9'd107: ReadData = 0;
9'd108: ReadData = 0;
9'd109: ReadData = 0;
9'd110: ReadData = 0;
9'd111: ReadData = 0;
9'd112: ReadData = 0;
9'd113: ReadData = 0;
9'd114: ReadData = 0;
9'd115: ReadData = 0;
9'd116: ReadData = 0;
9'd117: ReadData = 0;
9'd118: ReadData = 0;
9'd119: ReadData = 0;
9'd120: ReadData = 0;
9'd121: ReadData = 0;
9'd122: ReadData = 0;
9'd123: ReadData = 0;
9'd124: ReadData = 0;
9'd125: ReadData = 0;
9'd126: ReadData = 0;
9'd127: ReadData = 0;
9'd128: ReadData = 0;
9'd129: ReadData = 0;
9'd130: ReadData = 0;
9'd131: ReadData = 0;
9'd132: ReadData = 0;
9'd133: ReadData = 0;
9'd134: ReadData = 0;
9'd135: ReadData = 0;
9'd136: ReadData = 0;
9'd137: ReadData = 0;
9'd138: ReadData = 0;
9'd139: ReadData = 0;
9'd140: ReadData = 0;
9'd141: ReadData = 0;
9'd142: ReadData = 0;
9'd143: ReadData = 0;
9'd144: ReadData = 0;
9'd145: ReadData = 0;
9'd146: ReadData = 0;
9'd147: ReadData = 0;
9'd148: ReadData = 0;
9'd149: ReadData = 0;
9'd150: ReadData = 0;
9'd151: ReadData = 0;
9'd152: ReadData = 0;
9'd153: ReadData = 0;
9'd154: ReadData = 0;
9'd155: ReadData = 0;
9'd156: ReadData = 0;
9'd157: ReadData = 0;
9'd158: ReadData = 0;
9'd159: ReadData = 0;
9'd160: ReadData = 0;
9'd161: ReadData = 0;
9'd162: ReadData = 0;
9'd163: ReadData = 0;
9'd164: ReadData = 0;
9'd165: ReadData = 0;
9'd166: ReadData = 0;
9'd167: ReadData = 0;
9'd168: ReadData = 0;
9'd169: ReadData = 0;
9'd170: ReadData = 0;
9'd171: ReadData = 0;
9'd172: ReadData = 0;
9'd173: ReadData = 0;
9'd174: ReadData = 0;
9'd175: ReadData = 0;
9'd176: ReadData = 0;
9'd177: ReadData = 0;
9'd178: ReadData = 0;
9'd179: ReadData = 0;
9'd180: ReadData = 0;
9'd181: ReadData = 0;
9'd182: ReadData = 0;
9'd183: ReadData = 0;
9'd184: ReadData = 0;
9'd185: ReadData = 0;
9'd186: ReadData = 0;
9'd187: ReadData = 0;
9'd188: ReadData = 0;
9'd189: ReadData = 0;
9'd190: ReadData = 0;
9'd191: ReadData = 0;
9'd192: ReadData = 0;
9'd193: ReadData = 0;
9'd194: ReadData = 0;
9'd195: ReadData = 0;
9'd196: ReadData = 0;
9'd197: ReadData = 0;
9'd198: ReadData = 0;
9'd199: ReadData = 0;
9'd200: ReadData = 0;
9'd201: ReadData = 0;
9'd202: ReadData = 0;
9'd203: ReadData = 0;
9'd204: ReadData = 0;
9'd205: ReadData = 0;
9'd206: ReadData = 0;
9'd207: ReadData = 0;
9'd208: ReadData = 0;
9'd209: ReadData = 0;
9'd210: ReadData = 0;
9'd211: ReadData = 0;
9'd212: ReadData = 0;
9'd213: ReadData = 0;
9'd214: ReadData = 0;
9'd215: ReadData = 0;
9'd216: ReadData = 0;
9'd217: ReadData = 0;
9'd218: ReadData = 0;
9'd219: ReadData = 0;
9'd220: ReadData = 0;
9'd221: ReadData = 0;
9'd222: ReadData = 0;
9'd223: ReadData = 0;
9'd224: ReadData = 0;
9'd225: ReadData = 0;
9'd226: ReadData = 0;
9'd227: ReadData = 0;
9'd228: ReadData = 0;
9'd229: ReadData = 0;
9'd230: ReadData = 0;
9'd231: ReadData = 0;
9'd232: ReadData = 0;
9'd233: ReadData = 0;
9'd234: ReadData = 0;
9'd235: ReadData = 0;
9'd236: ReadData = 0;
9'd237: ReadData = 0;
9'd238: ReadData = 0;
9'd239: ReadData = 0;
9'd240: ReadData = 0;
9'd241: ReadData = 0;
9'd242: ReadData = 0;
9'd243: ReadData = 0;
9'd244: ReadData = 0;
9'd245: ReadData = 0;
9'd246: ReadData = 0;
9'd247: ReadData = 0;
9'd248: ReadData = 0;
9'd249: ReadData = 0;
9'd250: ReadData = 0;
9'd251: ReadData = 0;
9'd252: ReadData = 0;
9'd253: ReadData = 0;
9'd254: ReadData = 0;
9'd255: ReadData = 0;
9'd256: ReadData = 0;
9'd257: ReadData = 0;
9'd258: ReadData = 0;
9'd259: ReadData = 0;
9'd260: ReadData = 0;
9'd261: ReadData = 0;
9'd262: ReadData = 0;
9'd263: ReadData = 0;
9'd264: ReadData = 0;
9'd265: ReadData = 0;
9'd266: ReadData = 0;
9'd267: ReadData = 0;
9'd268: ReadData = 0;
9'd269: ReadData = 0;
9'd270: ReadData = 0;
9'd271: ReadData = 0;
9'd272: ReadData = 0;
9'd273: ReadData = 0;
9'd274: ReadData = 0;
9'd275: ReadData = 0;
9'd276: ReadData = 0;
9'd277: ReadData = 0;
9'd278: ReadData = 0;
9'd279: ReadData = 0;
9'd280: ReadData = 0;
9'd281: ReadData = 0;
9'd282: ReadData = 0;
9'd283: ReadData = 0;
9'd284: ReadData = 0;
9'd285: ReadData = 0;
9'd286: ReadData = 0;
9'd287: ReadData = 0;
9'd288: ReadData = 0;
9'd289: ReadData = 0;
9'd290: ReadData = 0;
9'd291: ReadData = 0;
9'd292: ReadData = 0;
9'd293: ReadData = 0;
9'd294: ReadData = 0;
9'd295: ReadData = 0;
9'd296: ReadData = 0;
9'd297: ReadData = 0;
9'd298: ReadData = 0;
9'd299: ReadData = 0;
9'd300: ReadData = 0;
9'd301: ReadData = 0;
9'd302: ReadData = 0;
9'd303: ReadData = 0;
9'd304: ReadData = 0;
9'd305: ReadData = 0;
9'd306: ReadData = 0;
9'd307: ReadData = 0;
9'd308: ReadData = 0;
9'd309: ReadData = 0;
9'd310: ReadData = 0;
9'd311: ReadData = 0;
9'd312: ReadData = 0;
9'd313: ReadData = 0;
9'd314: ReadData = 0;
9'd315: ReadData = 0;
9'd316: ReadData = 0;
9'd317: ReadData = 0;
9'd318: ReadData = 0;
9'd319: ReadData = 0;
9'd320: ReadData = 0;
9'd321: ReadData = 0;
9'd322: ReadData = 0;
9'd323: ReadData = 0;
9'd324: ReadData = 0;
9'd325: ReadData = 0;
9'd326: ReadData = 0;
9'd327: ReadData = 0;
9'd328: ReadData = 0;
9'd329: ReadData = 0;
9'd330: ReadData = 0;
9'd331: ReadData = 0;
9'd332: ReadData = 0;
9'd333: ReadData = 0;
9'd334: ReadData = 0;
9'd335: ReadData = 0;
9'd336: ReadData = 0;
9'd337: ReadData = 0;
9'd338: ReadData = 0;
9'd339: ReadData = 0;
9'd340: ReadData = 0;
9'd341: ReadData = 0;
9'd342: ReadData = 0;
9'd343: ReadData = 0;
9'd344: ReadData = 0;
9'd345: ReadData = 0;
9'd346: ReadData = 0;
9'd347: ReadData = 0;
9'd348: ReadData = 0;
9'd349: ReadData = 0;
9'd350: ReadData = 0;
9'd351: ReadData = 0;
9'd352: ReadData = 0;
9'd353: ReadData = 0;
9'd354: ReadData = 0;
9'd355: ReadData = 0;
9'd356: ReadData = 0;
9'd357: ReadData = 0;
9'd358: ReadData = 0;
9'd359: ReadData = 0;
9'd360: ReadData = 0;
9'd361: ReadData = 0;
9'd362: ReadData = 0;
9'd363: ReadData = 0;
9'd364: ReadData = 0;
9'd365: ReadData = 0;
9'd366: ReadData = 0;
9'd367: ReadData = 0;
9'd368: ReadData = 0;
9'd369: ReadData = 0;
9'd370: ReadData = 0;
9'd371: ReadData = 0;
9'd372: ReadData = 0;
9'd373: ReadData = 0;
9'd374: ReadData = 0;
9'd375: ReadData = 0;
9'd376: ReadData = 0;
9'd377: ReadData = 0;
9'd378: ReadData = 0;
9'd379: ReadData = 0;
9'd380: ReadData = 0;
9'd381: ReadData = 0;
9'd382: ReadData = 0;
9'd383: ReadData = 0;
9'd384: ReadData = 0;
9'd385: ReadData = 0;
9'd386: ReadData = 0;
9'd387: ReadData = 0;
9'd388: ReadData = 0;
9'd389: ReadData = 0;
9'd390: ReadData = 0;
9'd391: ReadData = 0;
9'd392: ReadData = 0;
9'd393: ReadData = 0;
9'd394: ReadData = 0;
9'd395: ReadData = 0;
9'd396: ReadData = 0;
9'd397: ReadData = 0;
9'd398: ReadData = 0;
9'd399: ReadData = 0;
9'd400: ReadData = 0;
9'd401: ReadData = 0;
9'd402: ReadData = 0;
9'd403: ReadData = 0;
9'd404: ReadData = 0;
9'd405: ReadData = 0;
9'd406: ReadData = 0;
9'd407: ReadData = 0;
9'd408: ReadData = 0;
9'd409: ReadData = 0;
9'd410: ReadData = 0;
9'd411: ReadData = 0;
9'd412: ReadData = 0;
9'd413: ReadData = 0;
9'd414: ReadData = 0;
9'd415: ReadData = 0;
9'd416: ReadData = 0;
9'd417: ReadData = 0;
9'd418: ReadData = 0;
9'd419: ReadData = 0;
9'd420: ReadData = 0;
9'd421: ReadData = 0;
9'd422: ReadData = 0;
9'd423: ReadData = 0;
9'd424: ReadData = 0;
9'd425: ReadData = 0;
9'd426: ReadData = 0;
9'd427: ReadData = 0;
9'd428: ReadData = 0;
9'd429: ReadData = 0;
9'd430: ReadData = 0;
9'd431: ReadData = 0;
9'd432: ReadData = 0;
9'd433: ReadData = 0;
9'd434: ReadData = 0;
9'd435: ReadData = 0;
9'd436: ReadData = 0;
9'd437: ReadData = 0;
9'd438: ReadData = 0;
9'd439: ReadData = 0;
9'd440: ReadData = 0;
9'd441: ReadData = 0;
9'd442: ReadData = 0;
9'd443: ReadData = 0;
9'd444: ReadData = 0;
9'd445: ReadData = 0;
9'd446: ReadData = 0;
9'd447: ReadData = 0;
9'd448: ReadData = 0;
9'd449: ReadData = 0;
9'd450: ReadData = 0;
9'd451: ReadData = 0;
9'd452: ReadData = 0;
9'd453: ReadData = 0;
9'd454: ReadData = 0;
9'd455: ReadData = 0;
9'd456: ReadData = 0;
9'd457: ReadData = 0;
9'd458: ReadData = 0;
9'd459: ReadData = 0;
9'd460: ReadData = 0;
9'd461: ReadData = 0;
9'd462: ReadData = 0;
9'd463: ReadData = 0;
9'd464: ReadData = 0;
9'd465: ReadData = 0;
9'd466: ReadData = 0;
9'd467: ReadData = 0;
9'd468: ReadData = 0;
9'd469: ReadData = 0;
9'd470: ReadData = 0;
9'd471: ReadData = 0;
9'd472: ReadData = 0;
9'd473: ReadData = 0;
9'd474: ReadData = 0;
9'd475: ReadData = 0;
9'd476: ReadData = 0;
9'd477: ReadData = 0;
9'd478: ReadData = 0;
9'd479: ReadData = 0;
9'd480: ReadData = 0;
9'd481: ReadData = 0;
9'd482: ReadData = 0;
9'd483: ReadData = 0;
9'd484: ReadData = 0;
9'd485: ReadData = 0;
9'd486: ReadData = 0;
9'd487: ReadData = 0;
9'd488: ReadData = 0;
9'd489: ReadData = 0;
9'd490: ReadData = 0;
9'd491: ReadData = 0;
9'd492: ReadData = 0;
9'd493: ReadData = 0;
9'd494: ReadData = 0;
9'd495: ReadData = 0;
9'd496: ReadData = 0;
9'd497: ReadData = 0;
9'd498: ReadData = 0;
9'd499: ReadData = 0;
9'd500: ReadData = 0;
9'd501: ReadData = 0;
9'd502: ReadData = 0;
9'd503: ReadData = 0;
9'd504: ReadData = 0;
9'd505: ReadData = 0;
9'd506: ReadData = 0;
9'd507: ReadData = 0;
9'd508: ReadData = 0;
9'd509: ReadData = 0;
9'd510: ReadData = 0;
9'd511: ReadData = 0;
endcase
end



endmodule
